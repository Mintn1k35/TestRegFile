library verilog;
use verilog.vl_types.all;
entity ifDut is
end ifDut;
